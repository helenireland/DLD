`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Digital Logic Design
// Engineer: Helen & Miguel
// 
// 7-segment display



// Create Date: 01/15/2021 06:40:11 PM
// Design Name: 
// Module Name: top_demo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top_demo
(
  // input
  input  logic [7:0] sw,
  input  logic [3:0] btn,
  input  logic       sysclk_125mhz,
  input  logic       rst,
  // output  
  output logic [7:0] led,
  output logic sseg_ca,
  output logic sseg_cb,
  output logic sseg_cc,
  output logic sseg_cd,
  output logic sseg_ce,
  output logic sseg_cf,
  output logic sseg_cg,
  output logic sseg_dp,
  output logic [3:0] sseg_an
);

  logic [16:0] CURRENT_COUNT;
  logic [16:0] NEXT_COUNT;
  logic        smol_clk;
  logic [3:0] sum;
  logic y;
  
  // Place TicTacToe instantiation here
  
  // 7-segment display
  segment_driver driver(
  .clk(smol_clk),
  .rst(btn[3]),
  .digit0(sw[3:0]),
  .digit1(sw[7:4]),
  .digit2(sum),
  .digit3(y),
  .decimals({1'b0, btn[2:0]}),
  .segment_cathodes({sseg_dp, sseg_cg, sseg_cf, sseg_ce, sseg_cd, sseg_cc, sseg_cb, sseg_ca}),
  .digit_anodes(sseg_an)
  );

// Register logic storing clock counts
  always@(posedge sysclk_125mhz)
  begin
    if(btn[3])
      CURRENT_COUNT = 17'h00000;
    else
      CURRENT_COUNT = NEXT_COUNT;
  end
  
  // Increment logic
  assign NEXT_COUNT = CURRENT_COUNT == 17'd100000 ? 17'h00000 : CURRENT_COUNT + 1;

  // Creation of smaller clock signal from counters
  assign smol_clk = CURRENT_COUNT == 17'd100000 ? 1'b1 : 1'b0;
  
 RCA dut(sw[3:0], sw[7:4], btn[0], y, sum);
 
endmodule
module RCA (input logic [3:0] a, b, input logic c, output logic y, output logic [3:0] sum);
  logic [2:0] cin;
  
  


  silly FA0 (a[0], b[0], c, cin[0], sum[0]); 
  silly FA1 (a[1], b[1], cin[0], cin[1], sum[1]);
  silly FA2 (a[2], b[2], cin[1], cin[2], sum[2]);
  silly FA3 (a[3], b[3], cin[2], y, sum[3]);
endmodule
module silly (input  logic a, b, c, output logic y, sum);
   
  assign sum = a ^ b ^ c;

  assign y = (a & b) | (a & c) | (b & c);
   
endmodule
